* inv.sp
*----------------------------------------------------------------------
* Parameters and models
*----------------------------------------------------------------------
.param SUPPLY=1.8
.lib 'rf018.l'  TT  
.temp 70

*----------------------------------------------------------------------
* Simulation netlist
*----------------------------------------------------------------------
Vgg vd gnd 'SUPPLY'
Vbb vb gnd -1

M1 vd vd gnd vb nch W=1000n L=180n

*----------------------------------------------------------------------
* Stimulus
*----------------------------------------------------------------------
.OP

.end